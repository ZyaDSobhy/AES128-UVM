
`include "sequence_item.sv"
 `include "driver.sv"
`include "monitor.sv"
  `include "sequence.sv"
 `include "sequencer.sv"
  `include "agent.sv"
`include "scoreboard.sv"
 `include "subscriber.sv"
`include "env.sv"
`include "test.sv"
